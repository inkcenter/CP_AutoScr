*.tran 0.1ps 1ns sweep monte=300
.tran 0.1ps 2ns

vX2_R/A X2_R/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX2_L/A X2_L/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX2_H/A X2_H/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX4_R/A X4_R/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX4_L/A X4_L/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX4_H/A X4_H/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX8_R/A X8_R/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX8_L/A X8_L/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX8_H/A X8_H/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX16_R/A X16_R/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX16_L/A X16_L/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX16_H/A X16_H/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX32_R/A X32_R/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX32_L/A X32_L/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

vX32_H/A X32_H/A 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

*sel=0
vXm4x1_R/S1 Xm4x1_R/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_R/S1 Xm4x2_R/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
*sel=1
vXm2x1_R/S0 Xm2x1_R/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm2x2_R/S0 Xm2x2_R/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x1_R/S0 Xm4x1_R/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x2_R/S0 Xm4x2_R/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
*A*=0
vXm2x1_R/A1 Xm2x1_R/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm2x2_R/A1 Xm2x2_R/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_R/A1 Xm4x1_R/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_R/A4 Xm4x1_R/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_R/A3 Xm4x1_R/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_R/A1 Xm4x2_R/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_R/A4 Xm4x2_R/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_R/A3 Xm4x2_R/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
*A2=1
vXm2x1_R/A2 Xm2x1_R/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm2x2_R/A2 Xm2x2_R/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x1_R/A2 Xm4x1_R/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x2_R/A2 Xm4x2_R/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

*LVT
vXm4x1_L/S1 Xm4x1_L/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_L/S1 Xm4x2_L/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)

vXm2x1_L/S0 Xm2x1_L/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm2x2_L/S0 Xm2x2_L/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x1_L/S0 Xm4x1_L/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x2_L/S0 Xm4x2_L/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)

vXm2x1_L/A1 Xm2x1_L/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm2x2_L/A1 Xm2x2_L/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_L/A1 Xm4x1_L/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_L/A4 Xm4x1_L/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_L/A3 Xm4x1_L/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_L/A1 Xm4x2_L/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_L/A4 Xm4x2_L/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_L/A3 Xm4x2_L/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)

vXm2x1_L/A2 Xm2x1_L/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm2x2_L/A2 Xm2x2_L/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x1_L/A2 Xm4x1_L/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x2_L/A2 Xm4x2_L/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

*HVT
vXm4x1_H/S1 Xm4x1_H/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_H/S1 Xm4x2_H/S1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)

vXm2x1_H/S0 Xm2x1_H/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm2x2_H/S0 Xm2x2_H/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x1_H/S0 Xm4x1_H/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)
vXm4x2_H/S0 Xm4x2_H/S0 0 PULSE (0 1.05 0.1ns 1ps 1ps 1ns 2ns)

vXm2x1_H/A1 Xm2x1_H/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm2x2_H/A1 Xm2x2_H/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_H/A1 Xm4x1_H/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_H/A4 Xm4x1_H/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x1_H/A3 Xm4x1_H/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_H/A1 Xm4x2_H/A1 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_H/A4 Xm4x2_H/A4 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)
vXm4x2_H/A3 Xm4x2_H/A3 0 PULSE (0 1.05 2ns 1ps 1ps 1ns 2ns)

vXm2x1_H/A2 Xm2x1_H/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm2x2_H/A2 Xm2x2_H/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x1_H/A2 Xm4x1_H/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)
vXm4x2_H/A2 Xm4x2_H/A2 0 pwl(0.0ns	0
+	0.50ns	0
+	0.50ns	0.0525
+	0.50ns	0.21
+	0.50ns	0.349146
+	0.50ns	0.470417
+	0.50ns	0.5775
+	0.50ns	0.673323
+	0.50ns	0.760208
+	0.50ns	0.84
+	0.50ns	0.914161
+	0.501ns	0.983854
+	0.501ns	1.05)

.measure tran delay_NBUFFX2_RVT
+ trig v(X2_R/A) val = 0.525 rise = 1
+ targ v(X2_R/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX2_LVT
+ trig v(X2_L/A) val = 0.525 rise = 1
+ targ v(X2_L/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX2_HVT
+ trig v(X2_H/A) val = 0.525 rise = 1
+ targ v(X2_H/Y) val = 0.525 rise = 1

.measure tran delay_NBUFFX4_RVT
+ trig v(X4_R/A) val = 0.525 rise = 1
+ targ v(X4_R/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX4_LVT
+ trig v(X4_L/A) val = 0.525 rise = 1
+ targ v(X4_L/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX4_HVT
+ trig v(X4_H/A) val = 0.525 rise = 1
+ targ v(X4_H/Y) val = 0.525 rise = 1

.measure tran delay_NBUFFX8_RVT
+ trig v(X8_R/A) val = 0.525 rise = 1
+ targ v(X8_R/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX8_LVT
+ trig v(X8_L/A) val = 0.525 rise = 1
+ targ v(X8_L/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX8_HVT
+ trig v(X8_H/A) val = 0.525 rise = 1
+ targ v(X8_H/Y) val = 0.525 rise = 1

.measure tran delay_NBUFFX16_RVT
+ trig v(X16_R/A) val = 0.525 rise = 1
+ targ v(X16_R/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX16_LVT
+ trig v(X16_L/A) val = 0.525 rise = 1
+ targ v(X16_L/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX16_HVT
+ trig v(X16_H/A) val = 0.525 rise = 1
+ targ v(X16_H/Y) val = 0.525 rise = 1

.measure tran delay_NBUFFX32_RVT
+ trig v(X32_R/A) val = 0.525 rise = 1
+ targ v(X32_R/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX32_LVT
+ trig v(X32_L/A) val = 0.525 rise = 1
+ targ v(X32_L/Y) val = 0.525 rise = 1
.measure tran delay_NBUFFX32_HVT
+ trig v(X32_H/A) val = 0.525 rise = 1
+ targ v(X32_H/Y) val = 0.525 rise = 1
*MUX_RVT
.measure tran delay_MUX21X1_RVT
+ trig v(Xm2x1_R/A2) val = 0.525 rise = 1
+ targ v(Xm2x1_R/Y) val = 0.525 rise = 1
.measure tran delay_MUX21X2_RVT
+ trig v(Xm2x2_R/A2) val = 0.525 rise = 1
+ targ v(Xm2x2_R/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X1_RVT
+ trig v(Xm4x1_R/A2) val = 0.525 rise = 1
+ targ v(Xm4x1_R/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X2_RVT
+ trig v(Xm4x2_R/A2) val = 0.525 rise = 1
+ targ v(Xm4x2_R/Y) val = 0.525 rise = 1
*MUX_LVT
.measure tran delay_MUX21X1_LVT
+ trig v(Xm2x1_L/A2) val = 0.525 rise = 1
+ targ v(Xm2x1_L/Y) val = 0.525 rise = 1
.measure tran delay_MUX21X2_LVT
+ trig v(Xm2x2_L/A2) val = 0.525 rise = 1
+ targ v(Xm2x2_L/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X1_LVT
+ trig v(Xm4x1_L/A2) val = 0.525 rise = 1
+ targ v(Xm4x1_L/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X2_LVT
+ trig v(Xm4x2_L/A2) val = 0.525 rise = 1
+ targ v(Xm4x2_L/Y) val = 0.525 rise = 1
*MUX_HVT
.measure tran delay_MUX21X1_HVT
+ trig v(Xm2x1_H/A2) val = 0.525 rise = 1
+ targ v(Xm2x1_H/Y) val = 0.525 rise = 1
.measure tran delay_MUX21X2_HVT
+ trig v(Xm2x2_H/A2) val = 0.525 rise = 1
+ targ v(Xm2x2_H/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X1_HVT
+ trig v(Xm4x1_H/A2) val = 0.525 rise = 1
+ targ v(Xm4x1_H/Y) val = 0.525 rise = 1
.measure tran delay_MUX41X2_HVT
+ trig v(Xm4x2_H/A2) val = 0.525 rise = 1
+ targ v(Xm4x2_H/Y) val = 0.525 rise = 1
