.tran 0.1ps 50ns

v000 000 0 PULSE ( 0 1.05 0.1ns 1ps 1ps 0.5ns 1ns )

